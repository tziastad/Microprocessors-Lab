library verilog;
use verilog.vl_types.all;
entity d1s4178tb2 is
end d1s4178tb2;
